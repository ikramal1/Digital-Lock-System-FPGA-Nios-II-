-- DigitalLock.vhd

-- Generated using ACDS version 13.0sp1 232 at 2026.01.22.00:32:32

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DigitalLock is
	port (
		clk_clk              : in  std_logic                     := '0';             --           clk.clk
		hex_external_export  : out std_logic_vector(27 downto 0);                    --  hex_external.export
		ledg_external_export : out std_logic_vector(7 downto 0);                     -- ledg_external.export
		ledr_external_export : out std_logic_vector(9 downto 0);                     -- ledr_external.export
		key_external_export  : in  std_logic_vector(3 downto 0)  := (others => '0'); --  key_external.export
		sw_external_export   : in  std_logic_vector(9 downto 0)  := (others => '0')  --   sw_external.export
	);
end entity DigitalLock;

architecture rtl of DigitalLock is
	component DigitalLock_CPU is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(14 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(14 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component DigitalLock_CPU;

	component DigitalLock_IN_RAM is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component DigitalLock_IN_RAM;

	component DigitalLock_JTAG_UART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component DigitalLock_JTAG_UART;

	component DigitalLock_HEX is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(27 downto 0)                     -- export
		);
	end component DigitalLock_HEX;

	component DigitalLock_LEDG is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component DigitalLock_LEDG;

	component DigitalLock_LEDR is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component DigitalLock_LEDR;

	component DigitalLock_KEY is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component DigitalLock_KEY;

	component DigitalLock_SW is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component DigitalLock_SW;

	component DigitalLock_TIMER is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component DigitalLock_TIMER;

	component DigitalLock_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component DigitalLock_sysid;

	component altera_merlin_master_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(89 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_agent;

	component altera_merlin_slave_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(14 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(89 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(90 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component altera_merlin_slave_agent;

	component altera_avalon_sc_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(90 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component altera_avalon_sc_fifo;

	component DigitalLock_addr_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(89 downto 0);                    -- data
			src_channel        : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component DigitalLock_addr_router;

	component DigitalLock_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(89 downto 0);                    -- data
			src_channel        : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component DigitalLock_addr_router_001;

	component DigitalLock_id_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(89 downto 0);                    -- data
			src_channel        : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component DigitalLock_id_router;

	component DigitalLock_id_router_002 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(89 downto 0);                    -- data
			src_channel        : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component DigitalLock_id_router_002;

	component DigitalLock_cmd_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(89 downto 0);                    -- data
			src0_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(89 downto 0);                    -- data
			src1_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component DigitalLock_cmd_xbar_demux;

	component DigitalLock_cmd_xbar_demux_001 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(89 downto 0);                    -- data
			src0_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(89 downto 0);                    -- data
			src1_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(89 downto 0);                    -- data
			src2_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic;                                        -- endofpacket
			src3_ready         : in  std_logic                     := 'X';             -- ready
			src3_valid         : out std_logic;                                        -- valid
			src3_data          : out std_logic_vector(89 downto 0);                    -- data
			src3_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src3_startofpacket : out std_logic;                                        -- startofpacket
			src3_endofpacket   : out std_logic;                                        -- endofpacket
			src4_ready         : in  std_logic                     := 'X';             -- ready
			src4_valid         : out std_logic;                                        -- valid
			src4_data          : out std_logic_vector(89 downto 0);                    -- data
			src4_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src4_startofpacket : out std_logic;                                        -- startofpacket
			src4_endofpacket   : out std_logic;                                        -- endofpacket
			src5_ready         : in  std_logic                     := 'X';             -- ready
			src5_valid         : out std_logic;                                        -- valid
			src5_data          : out std_logic_vector(89 downto 0);                    -- data
			src5_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src5_startofpacket : out std_logic;                                        -- startofpacket
			src5_endofpacket   : out std_logic;                                        -- endofpacket
			src6_ready         : in  std_logic                     := 'X';             -- ready
			src6_valid         : out std_logic;                                        -- valid
			src6_data          : out std_logic_vector(89 downto 0);                    -- data
			src6_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src6_startofpacket : out std_logic;                                        -- startofpacket
			src6_endofpacket   : out std_logic;                                        -- endofpacket
			src7_ready         : in  std_logic                     := 'X';             -- ready
			src7_valid         : out std_logic;                                        -- valid
			src7_data          : out std_logic_vector(89 downto 0);                    -- data
			src7_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src7_startofpacket : out std_logic;                                        -- startofpacket
			src7_endofpacket   : out std_logic;                                        -- endofpacket
			src8_ready         : in  std_logic                     := 'X';             -- ready
			src8_valid         : out std_logic;                                        -- valid
			src8_data          : out std_logic_vector(89 downto 0);                    -- data
			src8_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src8_startofpacket : out std_logic;                                        -- startofpacket
			src8_endofpacket   : out std_logic;                                        -- endofpacket
			src9_ready         : in  std_logic                     := 'X';             -- ready
			src9_valid         : out std_logic;                                        -- valid
			src9_data          : out std_logic_vector(89 downto 0);                    -- data
			src9_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src9_startofpacket : out std_logic;                                        -- startofpacket
			src9_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component DigitalLock_cmd_xbar_demux_001;

	component DigitalLock_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(89 downto 0);                    -- data
			src_channel         : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component DigitalLock_cmd_xbar_mux;

	component DigitalLock_rsp_xbar_demux_002 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(89 downto 0);                    -- data
			src0_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component DigitalLock_rsp_xbar_demux_002;

	component DigitalLock_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(89 downto 0);                    -- data
			src_channel         : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component DigitalLock_rsp_xbar_mux;

	component DigitalLock_rsp_xbar_mux_001 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(89 downto 0);                    -- data
			src_channel         : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                        -- ready
			sink3_valid         : in  std_logic                     := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready         : out std_logic;                                        -- ready
			sink4_valid         : in  std_logic                     := 'X';             -- valid
			sink4_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink4_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink4_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink5_ready         : out std_logic;                                        -- ready
			sink5_valid         : in  std_logic                     := 'X';             -- valid
			sink5_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink5_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink5_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink5_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink6_ready         : out std_logic;                                        -- ready
			sink6_valid         : in  std_logic                     := 'X';             -- valid
			sink6_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink6_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink6_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink6_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink7_ready         : out std_logic;                                        -- ready
			sink7_valid         : in  std_logic                     := 'X';             -- valid
			sink7_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink7_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink7_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink7_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink8_ready         : out std_logic;                                        -- ready
			sink8_valid         : in  std_logic                     := 'X';             -- valid
			sink8_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink8_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink8_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink8_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink9_ready         : out std_logic;                                        -- ready
			sink9_valid         : in  std_logic                     := 'X';             -- valid
			sink9_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink9_data          : in  std_logic_vector(89 downto 0) := (others => 'X'); -- data
			sink9_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink9_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component DigitalLock_rsp_xbar_mux_001;

	component DigitalLock_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component DigitalLock_irq_mapper;

	component digitallock_cpu_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(14 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component digitallock_cpu_instruction_master_translator;

	component digitallock_cpu_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(14 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component digitallock_cpu_data_master_translator;

	component digitallock_cpu_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component digitallock_cpu_jtag_debug_module_translator;

	component digitallock_in_ram_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(10 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component digitallock_in_ram_s1_translator;

	component digitallock_jtag_uart_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component digitallock_jtag_uart_avalon_jtag_slave_translator;

	component digitallock_hex_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component digitallock_hex_s1_translator;

	component digitallock_key_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component digitallock_key_s1_translator;

	component digitallock_timer_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component digitallock_timer_s1_translator;

	component digitallock_sysid_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component digitallock_sysid_control_slave_translator;

	component digitallock_rst_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component digitallock_rst_controller;

	component digitallock_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component digitallock_rst_controller_001;

	signal cpu_jtag_debug_module_reset_reset                                                                : std_logic;                     -- CPU:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	signal cpu_instruction_master_waitrequest                                                               : std_logic;                     -- CPU_instruction_master_translator:av_waitrequest -> CPU:i_waitrequest
	signal cpu_instruction_master_address                                                                   : std_logic_vector(14 downto 0); -- CPU:i_address -> CPU_instruction_master_translator:av_address
	signal cpu_instruction_master_read                                                                      : std_logic;                     -- CPU:i_read -> CPU_instruction_master_translator:av_read
	signal cpu_instruction_master_readdata                                                                  : std_logic_vector(31 downto 0); -- CPU_instruction_master_translator:av_readdata -> CPU:i_readdata
	signal cpu_data_master_waitrequest                                                                      : std_logic;                     -- CPU_data_master_translator:av_waitrequest -> CPU:d_waitrequest
	signal cpu_data_master_writedata                                                                        : std_logic_vector(31 downto 0); -- CPU:d_writedata -> CPU_data_master_translator:av_writedata
	signal cpu_data_master_address                                                                          : std_logic_vector(14 downto 0); -- CPU:d_address -> CPU_data_master_translator:av_address
	signal cpu_data_master_write                                                                            : std_logic;                     -- CPU:d_write -> CPU_data_master_translator:av_write
	signal cpu_data_master_read                                                                             : std_logic;                     -- CPU:d_read -> CPU_data_master_translator:av_read
	signal cpu_data_master_readdata                                                                         : std_logic_vector(31 downto 0); -- CPU_data_master_translator:av_readdata -> CPU:d_readdata
	signal cpu_data_master_debugaccess                                                                      : std_logic;                     -- CPU:jtag_debug_module_debugaccess_to_roms -> CPU_data_master_translator:av_debugaccess
	signal cpu_data_master_byteenable                                                                       : std_logic_vector(3 downto 0);  -- CPU:d_byteenable -> CPU_data_master_translator:av_byteenable
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                                 : std_logic;                     -- CPU:jtag_debug_module_waitrequest -> CPU_jtag_debug_module_translator:av_waitrequest
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata                                   : std_logic_vector(31 downto 0); -- CPU_jtag_debug_module_translator:av_writedata -> CPU:jtag_debug_module_writedata
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_address                                     : std_logic_vector(8 downto 0);  -- CPU_jtag_debug_module_translator:av_address -> CPU:jtag_debug_module_address
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_write                                       : std_logic;                     -- CPU_jtag_debug_module_translator:av_write -> CPU:jtag_debug_module_write
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_read                                        : std_logic;                     -- CPU_jtag_debug_module_translator:av_read -> CPU:jtag_debug_module_read
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata                                    : std_logic_vector(31 downto 0); -- CPU:jtag_debug_module_readdata -> CPU_jtag_debug_module_translator:av_readdata
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                                 : std_logic;                     -- CPU_jtag_debug_module_translator:av_debugaccess -> CPU:jtag_debug_module_debugaccess
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                                  : std_logic_vector(3 downto 0);  -- CPU_jtag_debug_module_translator:av_byteenable -> CPU:jtag_debug_module_byteenable
	signal in_ram_s1_translator_avalon_anti_slave_0_writedata                                               : std_logic_vector(31 downto 0); -- IN_RAM_s1_translator:av_writedata -> IN_RAM:writedata
	signal in_ram_s1_translator_avalon_anti_slave_0_address                                                 : std_logic_vector(10 downto 0); -- IN_RAM_s1_translator:av_address -> IN_RAM:address
	signal in_ram_s1_translator_avalon_anti_slave_0_chipselect                                              : std_logic;                     -- IN_RAM_s1_translator:av_chipselect -> IN_RAM:chipselect
	signal in_ram_s1_translator_avalon_anti_slave_0_clken                                                   : std_logic;                     -- IN_RAM_s1_translator:av_clken -> IN_RAM:clken
	signal in_ram_s1_translator_avalon_anti_slave_0_write                                                   : std_logic;                     -- IN_RAM_s1_translator:av_write -> IN_RAM:write
	signal in_ram_s1_translator_avalon_anti_slave_0_readdata                                                : std_logic_vector(31 downto 0); -- IN_RAM:readdata -> IN_RAM_s1_translator:av_readdata
	signal in_ram_s1_translator_avalon_anti_slave_0_byteenable                                              : std_logic_vector(3 downto 0);  -- IN_RAM_s1_translator:av_byteenable -> IN_RAM:byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                           : std_logic;                     -- JTAG_UART:av_waitrequest -> JTAG_UART_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0); -- JTAG_UART_avalon_jtag_slave_translator:av_writedata -> JTAG_UART:av_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address                               : std_logic_vector(0 downto 0);  -- JTAG_UART_avalon_jtag_slave_translator:av_address -> JTAG_UART:av_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                            : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator:av_chipselect -> JTAG_UART:av_chipselect
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                 : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator:av_write -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                  : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator:av_read -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0); -- JTAG_UART:av_readdata -> JTAG_UART_avalon_jtag_slave_translator:av_readdata
	signal hex_s1_translator_avalon_anti_slave_0_writedata                                                  : std_logic_vector(31 downto 0); -- HEX_s1_translator:av_writedata -> HEX:writedata
	signal hex_s1_translator_avalon_anti_slave_0_address                                                    : std_logic_vector(1 downto 0);  -- HEX_s1_translator:av_address -> HEX:address
	signal hex_s1_translator_avalon_anti_slave_0_chipselect                                                 : std_logic;                     -- HEX_s1_translator:av_chipselect -> HEX:chipselect
	signal hex_s1_translator_avalon_anti_slave_0_write                                                      : std_logic;                     -- HEX_s1_translator:av_write -> hex_s1_translator_avalon_anti_slave_0_write:in
	signal hex_s1_translator_avalon_anti_slave_0_readdata                                                   : std_logic_vector(31 downto 0); -- HEX:readdata -> HEX_s1_translator:av_readdata
	signal ledg_s1_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(31 downto 0); -- LEDG_s1_translator:av_writedata -> LEDG:writedata
	signal ledg_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(1 downto 0);  -- LEDG_s1_translator:av_address -> LEDG:address
	signal ledg_s1_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                     -- LEDG_s1_translator:av_chipselect -> LEDG:chipselect
	signal ledg_s1_translator_avalon_anti_slave_0_write                                                     : std_logic;                     -- LEDG_s1_translator:av_write -> ledg_s1_translator_avalon_anti_slave_0_write:in
	signal ledg_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(31 downto 0); -- LEDG:readdata -> LEDG_s1_translator:av_readdata
	signal ledr_s1_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(31 downto 0); -- LEDR_s1_translator:av_writedata -> LEDR:writedata
	signal ledr_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(1 downto 0);  -- LEDR_s1_translator:av_address -> LEDR:address
	signal ledr_s1_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                     -- LEDR_s1_translator:av_chipselect -> LEDR:chipselect
	signal ledr_s1_translator_avalon_anti_slave_0_write                                                     : std_logic;                     -- LEDR_s1_translator:av_write -> ledr_s1_translator_avalon_anti_slave_0_write:in
	signal ledr_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(31 downto 0); -- LEDR:readdata -> LEDR_s1_translator:av_readdata
	signal key_s1_translator_avalon_anti_slave_0_address                                                    : std_logic_vector(1 downto 0);  -- KEY_s1_translator:av_address -> KEY:address
	signal key_s1_translator_avalon_anti_slave_0_readdata                                                   : std_logic_vector(31 downto 0); -- KEY:readdata -> KEY_s1_translator:av_readdata
	signal sw_s1_translator_avalon_anti_slave_0_address                                                     : std_logic_vector(1 downto 0);  -- SW_s1_translator:av_address -> SW:address
	signal sw_s1_translator_avalon_anti_slave_0_readdata                                                    : std_logic_vector(31 downto 0); -- SW:readdata -> SW_s1_translator:av_readdata
	signal timer_s1_translator_avalon_anti_slave_0_writedata                                                : std_logic_vector(15 downto 0); -- TIMER_s1_translator:av_writedata -> TIMER:writedata
	signal timer_s1_translator_avalon_anti_slave_0_address                                                  : std_logic_vector(2 downto 0);  -- TIMER_s1_translator:av_address -> TIMER:address
	signal timer_s1_translator_avalon_anti_slave_0_chipselect                                               : std_logic;                     -- TIMER_s1_translator:av_chipselect -> TIMER:chipselect
	signal timer_s1_translator_avalon_anti_slave_0_write                                                    : std_logic;                     -- TIMER_s1_translator:av_write -> timer_s1_translator_avalon_anti_slave_0_write:in
	signal timer_s1_translator_avalon_anti_slave_0_readdata                                                 : std_logic_vector(15 downto 0); -- TIMER:readdata -> TIMER_s1_translator:av_readdata
	signal sysid_control_slave_translator_avalon_anti_slave_0_address                                       : std_logic_vector(0 downto 0);  -- sysid_control_slave_translator:av_address -> sysid:address
	signal sysid_control_slave_translator_avalon_anti_slave_0_readdata                                      : std_logic_vector(31 downto 0); -- sysid:readdata -> sysid_control_slave_translator:av_readdata
	signal cpu_instruction_master_translator_avalon_universal_master_0_waitrequest                          : std_logic;                     -- CPU_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_instruction_master_translator:uav_waitrequest
	signal cpu_instruction_master_translator_avalon_universal_master_0_burstcount                           : std_logic_vector(2 downto 0);  -- CPU_instruction_master_translator:uav_burstcount -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_instruction_master_translator_avalon_universal_master_0_writedata                            : std_logic_vector(31 downto 0); -- CPU_instruction_master_translator:uav_writedata -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_instruction_master_translator_avalon_universal_master_0_address                              : std_logic_vector(14 downto 0); -- CPU_instruction_master_translator:uav_address -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_instruction_master_translator_avalon_universal_master_0_lock                                 : std_logic;                     -- CPU_instruction_master_translator:uav_lock -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_instruction_master_translator_avalon_universal_master_0_write                                : std_logic;                     -- CPU_instruction_master_translator:uav_write -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_instruction_master_translator_avalon_universal_master_0_read                                 : std_logic;                     -- CPU_instruction_master_translator:uav_read -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdata                             : std_logic_vector(31 downto 0); -- CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_instruction_master_translator:uav_readdata
	signal cpu_instruction_master_translator_avalon_universal_master_0_debugaccess                          : std_logic;                     -- CPU_instruction_master_translator:uav_debugaccess -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_instruction_master_translator_avalon_universal_master_0_byteenable                           : std_logic_vector(3 downto 0);  -- CPU_instruction_master_translator:uav_byteenable -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid                        : std_logic;                     -- CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_instruction_master_translator:uav_readdatavalid
	signal cpu_data_master_translator_avalon_universal_master_0_waitrequest                                 : std_logic;                     -- CPU_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_data_master_translator:uav_waitrequest
	signal cpu_data_master_translator_avalon_universal_master_0_burstcount                                  : std_logic_vector(2 downto 0);  -- CPU_data_master_translator:uav_burstcount -> CPU_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_data_master_translator_avalon_universal_master_0_writedata                                   : std_logic_vector(31 downto 0); -- CPU_data_master_translator:uav_writedata -> CPU_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_data_master_translator_avalon_universal_master_0_address                                     : std_logic_vector(14 downto 0); -- CPU_data_master_translator:uav_address -> CPU_data_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_data_master_translator_avalon_universal_master_0_lock                                        : std_logic;                     -- CPU_data_master_translator:uav_lock -> CPU_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_data_master_translator_avalon_universal_master_0_write                                       : std_logic;                     -- CPU_data_master_translator:uav_write -> CPU_data_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_data_master_translator_avalon_universal_master_0_read                                        : std_logic;                     -- CPU_data_master_translator:uav_read -> CPU_data_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_data_master_translator_avalon_universal_master_0_readdata                                    : std_logic_vector(31 downto 0); -- CPU_data_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_data_master_translator:uav_readdata
	signal cpu_data_master_translator_avalon_universal_master_0_debugaccess                                 : std_logic;                     -- CPU_data_master_translator:uav_debugaccess -> CPU_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_data_master_translator_avalon_universal_master_0_byteenable                                  : std_logic_vector(3 downto 0);  -- CPU_data_master_translator:uav_byteenable -> CPU_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_data_master_translator_avalon_universal_master_0_readdatavalid                               : std_logic;                     -- CPU_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_data_master_translator:uav_readdatavalid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest                   : std_logic;                     -- CPU_jtag_debug_module_translator:uav_waitrequest -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount                    : std_logic_vector(2 downto 0);  -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> CPU_jtag_debug_module_translator:uav_burstcount
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata                     : std_logic_vector(31 downto 0); -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> CPU_jtag_debug_module_translator:uav_writedata
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                       : std_logic_vector(14 downto 0); -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> CPU_jtag_debug_module_translator:uav_address
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                         : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> CPU_jtag_debug_module_translator:uav_write
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                          : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> CPU_jtag_debug_module_translator:uav_lock
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                          : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> CPU_jtag_debug_module_translator:uav_read
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                      : std_logic_vector(31 downto 0); -- CPU_jtag_debug_module_translator:uav_readdata -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid                 : std_logic;                     -- CPU_jtag_debug_module_translator:uav_readdatavalid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess                   : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CPU_jtag_debug_module_translator:uav_debugaccess
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable                    : std_logic_vector(3 downto 0);  -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> CPU_jtag_debug_module_translator:uav_byteenable
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket            : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid                  : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket          : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data                   : std_logic_vector(90 downto 0); -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready                  : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket         : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid               : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket       : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                : std_logic_vector(90 downto 0); -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready               : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid             : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data              : std_logic_vector(33 downto 0); -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready             : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                               : std_logic;                     -- IN_RAM_s1_translator:uav_waitrequest -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                : std_logic_vector(2 downto 0);  -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> IN_RAM_s1_translator:uav_burstcount
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                 : std_logic_vector(31 downto 0); -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> IN_RAM_s1_translator:uav_writedata
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_m0_address                                   : std_logic_vector(14 downto 0); -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:m0_address -> IN_RAM_s1_translator:uav_address
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_m0_write                                     : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:m0_write -> IN_RAM_s1_translator:uav_write
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock                                      : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:m0_lock -> IN_RAM_s1_translator:uav_lock
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_m0_read                                      : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:m0_read -> IN_RAM_s1_translator:uav_read
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                  : std_logic_vector(31 downto 0); -- IN_RAM_s1_translator:uav_readdata -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                             : std_logic;                     -- IN_RAM_s1_translator:uav_readdatavalid -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                               : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> IN_RAM_s1_translator:uav_debugaccess
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                : std_logic_vector(3 downto 0);  -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> IN_RAM_s1_translator:uav_byteenable
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                        : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> IN_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                              : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> IN_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                      : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> IN_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data                               : std_logic_vector(90 downto 0); -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> IN_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                              : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                     : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                           : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                   : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                            : std_logic_vector(90 downto 0); -- IN_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                           : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> IN_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                         : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                          : std_logic_vector(33 downto 0); -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                         : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator:uav_waitrequest -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);  -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> JTAG_UART_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0); -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> JTAG_UART_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(14 downto 0); -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> JTAG_UART_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> JTAG_UART_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> JTAG_UART_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> JTAG_UART_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0); -- JTAG_UART_avalon_jtag_slave_translator:uav_readdata -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator:uav_readdatavalid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> JTAG_UART_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);  -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> JTAG_UART_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(90 downto 0); -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(90 downto 0); -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0); -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal hex_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                     -- HEX_s1_translator:uav_waitrequest -> HEX_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal hex_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(2 downto 0);  -- HEX_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> HEX_s1_translator:uav_burstcount
	signal hex_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(31 downto 0); -- HEX_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> HEX_s1_translator:uav_writedata
	signal hex_s1_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(14 downto 0); -- HEX_s1_translator_avalon_universal_slave_0_agent:m0_address -> HEX_s1_translator:uav_address
	signal hex_s1_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:m0_write -> HEX_s1_translator:uav_write
	signal hex_s1_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:m0_lock -> HEX_s1_translator:uav_lock
	signal hex_s1_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:m0_read -> HEX_s1_translator:uav_read
	signal hex_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(31 downto 0); -- HEX_s1_translator:uav_readdata -> HEX_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal hex_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                     -- HEX_s1_translator:uav_readdatavalid -> HEX_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal hex_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> HEX_s1_translator:uav_debugaccess
	signal hex_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(3 downto 0);  -- HEX_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> HEX_s1_translator:uav_byteenable
	signal hex_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> HEX_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal hex_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> HEX_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal hex_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> HEX_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal hex_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(90 downto 0); -- HEX_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> HEX_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal hex_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> HEX_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> HEX_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> HEX_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> HEX_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(90 downto 0); -- HEX_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> HEX_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> HEX_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal hex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> HEX_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal hex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(33 downto 0); -- HEX_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> HEX_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal hex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> HEX_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                     -- LEDG_s1_translator:uav_waitrequest -> LEDG_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);  -- LEDG_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LEDG_s1_translator:uav_burstcount
	signal ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0); -- LEDG_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LEDG_s1_translator:uav_writedata
	signal ledg_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(14 downto 0); -- LEDG_s1_translator_avalon_universal_slave_0_agent:m0_address -> LEDG_s1_translator:uav_address
	signal ledg_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:m0_write -> LEDG_s1_translator:uav_write
	signal ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LEDG_s1_translator:uav_lock
	signal ledg_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:m0_read -> LEDG_s1_translator:uav_read
	signal ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0); -- LEDG_s1_translator:uav_readdata -> LEDG_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                     -- LEDG_s1_translator:uav_readdatavalid -> LEDG_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LEDG_s1_translator:uav_debugaccess
	signal ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);  -- LEDG_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LEDG_s1_translator:uav_byteenable
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(90 downto 0); -- LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(90 downto 0); -- LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0); -- LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                     -- LEDR_s1_translator:uav_waitrequest -> LEDR_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);  -- LEDR_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LEDR_s1_translator:uav_burstcount
	signal ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0); -- LEDR_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LEDR_s1_translator:uav_writedata
	signal ledr_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(14 downto 0); -- LEDR_s1_translator_avalon_universal_slave_0_agent:m0_address -> LEDR_s1_translator:uav_address
	signal ledr_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:m0_write -> LEDR_s1_translator:uav_write
	signal ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LEDR_s1_translator:uav_lock
	signal ledr_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:m0_read -> LEDR_s1_translator:uav_read
	signal ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0); -- LEDR_s1_translator:uav_readdata -> LEDR_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                     -- LEDR_s1_translator:uav_readdatavalid -> LEDR_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LEDR_s1_translator:uav_debugaccess
	signal ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);  -- LEDR_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LEDR_s1_translator:uav_byteenable
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(90 downto 0); -- LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(90 downto 0); -- LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0); -- LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                     -- KEY_s1_translator:uav_waitrequest -> KEY_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(2 downto 0);  -- KEY_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> KEY_s1_translator:uav_burstcount
	signal key_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(31 downto 0); -- KEY_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> KEY_s1_translator:uav_writedata
	signal key_s1_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(14 downto 0); -- KEY_s1_translator_avalon_universal_slave_0_agent:m0_address -> KEY_s1_translator:uav_address
	signal key_s1_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:m0_write -> KEY_s1_translator:uav_write
	signal key_s1_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:m0_lock -> KEY_s1_translator:uav_lock
	signal key_s1_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:m0_read -> KEY_s1_translator:uav_read
	signal key_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(31 downto 0); -- KEY_s1_translator:uav_readdata -> KEY_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                     -- KEY_s1_translator:uav_readdatavalid -> KEY_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> KEY_s1_translator:uav_debugaccess
	signal key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(3 downto 0);  -- KEY_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> KEY_s1_translator:uav_byteenable
	signal key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> KEY_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> KEY_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> KEY_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal key_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(90 downto 0); -- KEY_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> KEY_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> KEY_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> KEY_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> KEY_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> KEY_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(90 downto 0); -- KEY_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> KEY_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> KEY_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> KEY_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(33 downto 0); -- KEY_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> KEY_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> KEY_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                   : std_logic;                     -- SW_s1_translator:uav_waitrequest -> SW_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                    : std_logic_vector(2 downto 0);  -- SW_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SW_s1_translator:uav_burstcount
	signal sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                     : std_logic_vector(31 downto 0); -- SW_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SW_s1_translator:uav_writedata
	signal sw_s1_translator_avalon_universal_slave_0_agent_m0_address                                       : std_logic_vector(14 downto 0); -- SW_s1_translator_avalon_universal_slave_0_agent:m0_address -> SW_s1_translator:uav_address
	signal sw_s1_translator_avalon_universal_slave_0_agent_m0_write                                         : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:m0_write -> SW_s1_translator:uav_write
	signal sw_s1_translator_avalon_universal_slave_0_agent_m0_lock                                          : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SW_s1_translator:uav_lock
	signal sw_s1_translator_avalon_universal_slave_0_agent_m0_read                                          : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:m0_read -> SW_s1_translator:uav_read
	signal sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                      : std_logic_vector(31 downto 0); -- SW_s1_translator:uav_readdata -> SW_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                 : std_logic;                     -- SW_s1_translator:uav_readdatavalid -> SW_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                   : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SW_s1_translator:uav_debugaccess
	signal sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                    : std_logic_vector(3 downto 0);  -- SW_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SW_s1_translator:uav_byteenable
	signal sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                            : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                  : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                          : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                   : std_logic_vector(90 downto 0); -- SW_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                  : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SW_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                         : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                               : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                       : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                : std_logic_vector(90 downto 0); -- SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                               : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                             : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                              : std_logic_vector(33 downto 0); -- SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                             : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                : std_logic;                     -- TIMER_s1_translator:uav_waitrequest -> TIMER_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                 : std_logic_vector(2 downto 0);  -- TIMER_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> TIMER_s1_translator:uav_burstcount
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                  : std_logic_vector(31 downto 0); -- TIMER_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> TIMER_s1_translator:uav_writedata
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_address                                    : std_logic_vector(14 downto 0); -- TIMER_s1_translator_avalon_universal_slave_0_agent:m0_address -> TIMER_s1_translator:uav_address
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_write                                      : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:m0_write -> TIMER_s1_translator:uav_write
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_lock                                       : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:m0_lock -> TIMER_s1_translator:uav_lock
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_read                                       : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:m0_read -> TIMER_s1_translator:uav_read
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                   : std_logic_vector(31 downto 0); -- TIMER_s1_translator:uav_readdata -> TIMER_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                              : std_logic;                     -- TIMER_s1_translator:uav_readdatavalid -> TIMER_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> TIMER_s1_translator:uav_debugaccess
	signal timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                 : std_logic_vector(3 downto 0);  -- TIMER_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> TIMER_s1_translator:uav_byteenable
	signal timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                         : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                               : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                       : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                : std_logic_vector(90 downto 0); -- TIMER_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                               : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> TIMER_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                      : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> TIMER_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                            : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> TIMER_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                    : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> TIMER_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                             : std_logic_vector(90 downto 0); -- TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> TIMER_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                            : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                          : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> TIMER_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                           : std_logic_vector(33 downto 0); -- TIMER_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> TIMER_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                          : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> TIMER_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                     : std_logic;                     -- sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                      : std_logic_vector(2 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                       : std_logic_vector(31 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address                         : std_logic_vector(14 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write                           : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                            : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read                            : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                        : std_logic_vector(31 downto 0); -- sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                   : std_logic;                     -- sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                     : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                      : std_logic_vector(3 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket              : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                    : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket            : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                     : std_logic_vector(90 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                    : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket           : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                 : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket         : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                  : std_logic_vector(90 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                 : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid               : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                : std_logic_vector(33 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready               : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket                 : std_logic;                     -- CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                       : std_logic;                     -- CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket               : std_logic;                     -- CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data                        : std_logic_vector(89 downto 0); -- CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                       : std_logic;                     -- addr_router:sink_ready -> CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                        : std_logic;                     -- CPU_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid                              : std_logic;                     -- CPU_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                      : std_logic;                     -- CPU_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_data                               : std_logic_vector(89 downto 0); -- CPU_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready                              : std_logic;                     -- addr_router_001:sink_ready -> CPU_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket                   : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                         : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket                 : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                          : std_logic_vector(89 downto 0); -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                         : std_logic;                     -- id_router:sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                               : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid                                     : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                             : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rp_data                                      : std_logic_vector(89 downto 0); -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal in_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready                                     : std_logic;                     -- id_router_001:sink_ready -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(89 downto 0); -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                     -- id_router_002:sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal hex_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal hex_s1_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal hex_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal hex_s1_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(89 downto 0); -- HEX_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal hex_s1_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                     -- id_router_003:sink_ready -> HEX_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(89 downto 0); -- LEDG_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                     -- id_router_004:sink_ready -> LEDG_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(89 downto 0); -- LEDR_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                     -- id_router_005:sink_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal key_s1_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal key_s1_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(89 downto 0); -- KEY_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal key_s1_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                     -- id_router_006:sink_ready -> KEY_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                   : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal sw_s1_translator_avalon_universal_slave_0_agent_rp_valid                                         : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                 : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal sw_s1_translator_avalon_universal_slave_0_agent_rp_data                                          : std_logic_vector(89 downto 0); -- SW_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal sw_s1_translator_avalon_universal_slave_0_agent_rp_ready                                         : std_logic;                     -- id_router_007:sink_ready -> SW_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal timer_s1_translator_avalon_universal_slave_0_agent_rp_valid                                      : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                              : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal timer_s1_translator_avalon_universal_slave_0_agent_rp_data                                       : std_logic_vector(89 downto 0); -- TIMER_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal timer_s1_translator_avalon_universal_slave_0_agent_rp_ready                                      : std_logic;                     -- id_router_008:sink_ready -> TIMER_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                     : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                           : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                   : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data                            : std_logic_vector(89 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                           : std_logic;                     -- id_router_009:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal rst_controller_reset_out_reset                                                                   : std_logic;                     -- rst_controller:reset_out -> [CPU_data_master_translator:reset, CPU_data_master_translator_avalon_universal_master_0_agent:reset, CPU_instruction_master_translator:reset, CPU_instruction_master_translator_avalon_universal_master_0_agent:reset, CPU_jtag_debug_module_translator:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, id_router:reset, irq_mapper:reset, rsp_xbar_demux:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                                                               : std_logic;                     -- rst_controller_001:reset_out -> [HEX_s1_translator:reset, HEX_s1_translator_avalon_universal_slave_0_agent:reset, HEX_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, IN_RAM:reset, IN_RAM_s1_translator:reset, IN_RAM_s1_translator_avalon_universal_slave_0_agent:reset, IN_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, JTAG_UART_avalon_jtag_slave_translator:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, KEY_s1_translator:reset, KEY_s1_translator_avalon_universal_slave_0_agent:reset, KEY_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LEDG_s1_translator:reset, LEDG_s1_translator_avalon_universal_slave_0_agent:reset, LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LEDR_s1_translator:reset, LEDR_s1_translator_avalon_universal_slave_0_agent:reset, LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SW_s1_translator:reset, SW_s1_translator_avalon_universal_slave_0_agent:reset, SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, TIMER_s1_translator:reset, TIMER_s1_translator_avalon_universal_slave_0_agent:reset, TIMER_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_001:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rst_controller_001_reset_out_reset:in, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	signal rst_controller_001_reset_out_reset_req                                                           : std_logic;                     -- rst_controller_001:reset_req -> IN_RAM:reset_req
	signal cmd_xbar_demux_src0_endofpacket                                                                  : std_logic;                     -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                        : std_logic;                     -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                : std_logic;                     -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                         : std_logic_vector(89 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                      : std_logic_vector(9 downto 0);  -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                        : std_logic;                     -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                  : std_logic;                     -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                        : std_logic;                     -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                : std_logic;                     -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                         : std_logic_vector(89 downto 0); -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                      : std_logic_vector(9 downto 0);  -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                        : std_logic;                     -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                     : std_logic_vector(89 downto 0); -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                  : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                    : std_logic;                     -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                     : std_logic_vector(89 downto 0); -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                  : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                    : std_logic;                     -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src2_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src2_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src2_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                     : std_logic_vector(89 downto 0); -- cmd_xbar_demux_001:src2_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src2_channel                                                                  : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src2_channel -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src3_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src3_endofpacket -> HEX_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src3_valid -> HEX_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src3_startofpacket -> HEX_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                     : std_logic_vector(89 downto 0); -- cmd_xbar_demux_001:src3_data -> HEX_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src3_channel                                                                  : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src3_channel -> HEX_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src4_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src4_endofpacket -> LEDG_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src4_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src4_valid -> LEDG_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src4_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src4_startofpacket -> LEDG_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src4_data                                                                     : std_logic_vector(89 downto 0); -- cmd_xbar_demux_001:src4_data -> LEDG_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src4_channel                                                                  : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src4_channel -> LEDG_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src5_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src5_endofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src5_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src5_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src5_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src5_startofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src5_data                                                                     : std_logic_vector(89 downto 0); -- cmd_xbar_demux_001:src5_data -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src5_channel                                                                  : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src5_channel -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src6_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src6_endofpacket -> KEY_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src6_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src6_valid -> KEY_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src6_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src6_startofpacket -> KEY_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src6_data                                                                     : std_logic_vector(89 downto 0); -- cmd_xbar_demux_001:src6_data -> KEY_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src6_channel                                                                  : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src6_channel -> KEY_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src7_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src7_endofpacket -> SW_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src7_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src7_valid -> SW_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src7_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src7_startofpacket -> SW_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src7_data                                                                     : std_logic_vector(89 downto 0); -- cmd_xbar_demux_001:src7_data -> SW_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src7_channel                                                                  : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src7_channel -> SW_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src8_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src8_endofpacket -> TIMER_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src8_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src8_valid -> TIMER_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src8_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src8_startofpacket -> TIMER_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src8_data                                                                     : std_logic_vector(89 downto 0); -- cmd_xbar_demux_001:src8_data -> TIMER_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src8_channel                                                                  : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src8_channel -> TIMER_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src9_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src9_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src9_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src9_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src9_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src9_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src9_data                                                                     : std_logic_vector(89 downto 0); -- cmd_xbar_demux_001:src9_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src9_channel                                                                  : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src9_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal rsp_xbar_demux_src0_endofpacket                                                                  : std_logic;                     -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                        : std_logic;                     -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                : std_logic;                     -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                         : std_logic_vector(89 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                      : std_logic_vector(9 downto 0);  -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                        : std_logic;                     -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                  : std_logic;                     -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                        : std_logic;                     -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                : std_logic;                     -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                         : std_logic_vector(89 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                      : std_logic_vector(9 downto 0);  -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                        : std_logic;                     -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                              : std_logic;                     -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                    : std_logic;                     -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                            : std_logic;                     -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                     : std_logic_vector(89 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                  : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                    : std_logic;                     -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                              : std_logic;                     -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                    : std_logic;                     -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                            : std_logic;                     -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                     : std_logic_vector(89 downto 0); -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                  : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                    : std_logic;                     -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                              : std_logic;                     -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                    : std_logic;                     -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                            : std_logic;                     -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                     : std_logic_vector(89 downto 0); -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                  : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                    : std_logic;                     -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                              : std_logic;                     -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                    : std_logic;                     -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                            : std_logic;                     -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                     : std_logic_vector(89 downto 0); -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                  : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                    : std_logic;                     -- rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                              : std_logic;                     -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                    : std_logic;                     -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                            : std_logic;                     -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                     : std_logic_vector(89 downto 0); -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                  : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                    : std_logic;                     -- rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                              : std_logic;                     -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                    : std_logic;                     -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                            : std_logic;                     -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                     : std_logic_vector(89 downto 0); -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                                  : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                    : std_logic;                     -- rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                              : std_logic;                     -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                    : std_logic;                     -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                            : std_logic;                     -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                     : std_logic_vector(89 downto 0); -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                                  : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                    : std_logic;                     -- rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                              : std_logic;                     -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                    : std_logic;                     -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                            : std_logic;                     -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                     : std_logic_vector(89 downto 0); -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	signal rsp_xbar_demux_007_src0_channel                                                                  : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	signal rsp_xbar_demux_007_src0_ready                                                                    : std_logic;                     -- rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                              : std_logic;                     -- rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                    : std_logic;                     -- rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                            : std_logic;                     -- rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                     : std_logic_vector(89 downto 0); -- rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	signal rsp_xbar_demux_008_src0_channel                                                                  : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	signal rsp_xbar_demux_008_src0_ready                                                                    : std_logic;                     -- rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                              : std_logic;                     -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                    : std_logic;                     -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                            : std_logic;                     -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                     : std_logic_vector(89 downto 0); -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	signal rsp_xbar_demux_009_src0_channel                                                                  : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	signal rsp_xbar_demux_009_src0_ready                                                                    : std_logic;                     -- rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	signal addr_router_src_endofpacket                                                                      : std_logic;                     -- addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal addr_router_src_valid                                                                            : std_logic;                     -- addr_router:src_valid -> cmd_xbar_demux:sink_valid
	signal addr_router_src_startofpacket                                                                    : std_logic;                     -- addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal addr_router_src_data                                                                             : std_logic_vector(89 downto 0); -- addr_router:src_data -> cmd_xbar_demux:sink_data
	signal addr_router_src_channel                                                                          : std_logic_vector(9 downto 0);  -- addr_router:src_channel -> cmd_xbar_demux:sink_channel
	signal addr_router_src_ready                                                                            : std_logic;                     -- cmd_xbar_demux:sink_ready -> addr_router:src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                     : std_logic;                     -- rsp_xbar_mux:src_endofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_src_valid                                                                           : std_logic;                     -- rsp_xbar_mux:src_valid -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_src_startofpacket                                                                   : std_logic;                     -- rsp_xbar_mux:src_startofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_src_data                                                                            : std_logic_vector(89 downto 0); -- rsp_xbar_mux:src_data -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_src_channel                                                                         : std_logic_vector(9 downto 0);  -- rsp_xbar_mux:src_channel -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_src_ready                                                                           : std_logic;                     -- CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	signal addr_router_001_src_endofpacket                                                                  : std_logic;                     -- addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal addr_router_001_src_valid                                                                        : std_logic;                     -- addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	signal addr_router_001_src_startofpacket                                                                : std_logic;                     -- addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal addr_router_001_src_data                                                                         : std_logic_vector(89 downto 0); -- addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	signal addr_router_001_src_channel                                                                      : std_logic_vector(9 downto 0);  -- addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	signal addr_router_001_src_ready                                                                        : std_logic;                     -- cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                 : std_logic;                     -- rsp_xbar_mux_001:src_endofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                       : std_logic;                     -- rsp_xbar_mux_001:src_valid -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                               : std_logic;                     -- rsp_xbar_mux_001:src_startofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                        : std_logic_vector(89 downto 0); -- rsp_xbar_mux_001:src_data -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_001_src_channel                                                                     : std_logic_vector(9 downto 0);  -- rsp_xbar_mux_001:src_channel -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_001_src_ready                                                                       : std_logic;                     -- CPU_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                     : std_logic;                     -- cmd_xbar_mux:src_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                           : std_logic;                     -- cmd_xbar_mux:src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                   : std_logic;                     -- cmd_xbar_mux:src_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                            : std_logic_vector(89 downto 0); -- cmd_xbar_mux:src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                         : std_logic_vector(9 downto 0);  -- cmd_xbar_mux:src_channel -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                           : std_logic;                     -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                        : std_logic;                     -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                              : std_logic;                     -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                      : std_logic;                     -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                               : std_logic_vector(89 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                            : std_logic_vector(9 downto 0);  -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                              : std_logic;                     -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                 : std_logic;                     -- cmd_xbar_mux_001:src_endofpacket -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                       : std_logic;                     -- cmd_xbar_mux_001:src_valid -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                               : std_logic;                     -- cmd_xbar_mux_001:src_startofpacket -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                        : std_logic_vector(89 downto 0); -- cmd_xbar_mux_001:src_data -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_001_src_channel                                                                     : std_logic_vector(9 downto 0);  -- cmd_xbar_mux_001:src_channel -> IN_RAM_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_001_src_ready                                                                       : std_logic;                     -- IN_RAM_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                                    : std_logic;                     -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                          : std_logic;                     -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                  : std_logic;                     -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                           : std_logic_vector(89 downto 0); -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                        : std_logic_vector(9 downto 0);  -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                          : std_logic;                     -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_demux_001_src2_ready                                                                    : std_logic;                     -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	signal id_router_002_src_endofpacket                                                                    : std_logic;                     -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                          : std_logic;                     -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                  : std_logic;                     -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                           : std_logic_vector(89 downto 0); -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                        : std_logic_vector(9 downto 0);  -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                          : std_logic;                     -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal cmd_xbar_demux_001_src3_ready                                                                    : std_logic;                     -- HEX_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	signal id_router_003_src_endofpacket                                                                    : std_logic;                     -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                          : std_logic;                     -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                  : std_logic;                     -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                           : std_logic_vector(89 downto 0); -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                        : std_logic_vector(9 downto 0);  -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                          : std_logic;                     -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_demux_001_src4_ready                                                                    : std_logic;                     -- LEDG_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	signal id_router_004_src_endofpacket                                                                    : std_logic;                     -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                          : std_logic;                     -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                  : std_logic;                     -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                           : std_logic_vector(89 downto 0); -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                        : std_logic_vector(9 downto 0);  -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                          : std_logic;                     -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_demux_001_src5_ready                                                                    : std_logic;                     -- LEDR_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	signal id_router_005_src_endofpacket                                                                    : std_logic;                     -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                          : std_logic;                     -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                  : std_logic;                     -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                           : std_logic_vector(89 downto 0); -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                        : std_logic_vector(9 downto 0);  -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                          : std_logic;                     -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_demux_001_src6_ready                                                                    : std_logic;                     -- KEY_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	signal id_router_006_src_endofpacket                                                                    : std_logic;                     -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                          : std_logic;                     -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                  : std_logic;                     -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                           : std_logic_vector(89 downto 0); -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                        : std_logic_vector(9 downto 0);  -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                          : std_logic;                     -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_demux_001_src7_ready                                                                    : std_logic;                     -- SW_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	signal id_router_007_src_endofpacket                                                                    : std_logic;                     -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                          : std_logic;                     -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                  : std_logic;                     -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                           : std_logic_vector(89 downto 0); -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                        : std_logic_vector(9 downto 0);  -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                          : std_logic;                     -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_demux_001_src8_ready                                                                    : std_logic;                     -- TIMER_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	signal id_router_008_src_endofpacket                                                                    : std_logic;                     -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                          : std_logic;                     -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                  : std_logic;                     -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                           : std_logic_vector(89 downto 0); -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                        : std_logic_vector(9 downto 0);  -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                          : std_logic;                     -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_demux_001_src9_ready                                                                    : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	signal id_router_009_src_endofpacket                                                                    : std_logic;                     -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                          : std_logic;                     -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                  : std_logic;                     -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                           : std_logic_vector(89 downto 0); -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                        : std_logic_vector(9 downto 0);  -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                          : std_logic;                     -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal irq_mapper_receiver0_irq                                                                         : std_logic;                     -- JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                         : std_logic;                     -- TIMER:irq -> irq_mapper:receiver1_irq
	signal cpu_d_irq_irq                                                                                    : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> CPU:d_irq
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                       : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> JTAG_UART:av_write_n
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                        : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> JTAG_UART:av_read_n
	signal hex_s1_translator_avalon_anti_slave_0_write_ports_inv                                            : std_logic;                     -- hex_s1_translator_avalon_anti_slave_0_write:inv -> HEX:write_n
	signal ledg_s1_translator_avalon_anti_slave_0_write_ports_inv                                           : std_logic;                     -- ledg_s1_translator_avalon_anti_slave_0_write:inv -> LEDG:write_n
	signal ledr_s1_translator_avalon_anti_slave_0_write_ports_inv                                           : std_logic;                     -- ledr_s1_translator_avalon_anti_slave_0_write:inv -> LEDR:write_n
	signal timer_s1_translator_avalon_anti_slave_0_write_ports_inv                                          : std_logic;                     -- timer_s1_translator_avalon_anti_slave_0_write:inv -> TIMER:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                         : std_logic;                     -- rst_controller_reset_out_reset:inv -> CPU:reset_n
	signal rst_controller_001_reset_out_reset_ports_inv                                                     : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [HEX:reset_n, JTAG_UART:rst_n, KEY:reset_n, LEDG:reset_n, LEDR:reset_n, SW:reset_n, TIMER:reset_n, sysid:reset_n]

begin

	cpu : component DigitalLock_CPU
		port map (
			clk                                   => clk_clk,                                                          --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                         --                   reset_n.reset_n
			d_address                             => cpu_data_master_address,                                          --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                                       --                          .byteenable
			d_read                                => cpu_data_master_read,                                             --                          .read
			d_readdata                            => cpu_data_master_readdata,                                         --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                                      --                          .waitrequest
			d_write                               => cpu_data_master_write,                                            --                          .write
			d_writedata                           => cpu_data_master_writedata,                                        --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                                      --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                                   --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                                      --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                                  --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                               --                          .waitrequest
			d_irq                                 => cpu_d_irq_irq,                                                    --                     d_irq.irq
			jtag_debug_module_resetrequest        => cpu_jtag_debug_module_reset_reset,                                --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                          .read
			jtag_debug_module_readdata            => cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                          .write
			jtag_debug_module_writedata           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                          .writedata
			no_ci_readra                          => open                                                              -- custom_instruction_master.readra
		);

	in_ram : component DigitalLock_IN_RAM
		port map (
			clk        => clk_clk,                                             --   clk1.clk
			address    => in_ram_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			clken      => in_ram_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			chipselect => in_ram_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			write      => in_ram_s1_translator_avalon_anti_slave_0_write,      --       .write
			readdata   => in_ram_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			writedata  => in_ram_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => in_ram_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,                  -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req               --       .reset_req
		);

	jtag_uart : component DigitalLock_JTAG_UART
		port map (
			clk            => clk_clk,                                                                    --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                               --             reset.reset_n
			av_chipselect  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                                    --               irq.irq
		);

	hex : component DigitalLock_HEX
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => hex_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => hex_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => hex_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => hex_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => hex_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => hex_external_export                                    -- external_connection.export
		);

	ledg : component DigitalLock_LEDG
		port map (
			clk        => clk_clk,                                                --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => ledg_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => ledg_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => ledg_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => ledg_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => ledg_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => ledg_external_export                                    -- external_connection.export
		);

	ledr : component DigitalLock_LEDR
		port map (
			clk        => clk_clk,                                                --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => ledr_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => ledr_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => ledr_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => ledr_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => ledr_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => ledr_external_export                                    -- external_connection.export
		);

	key : component DigitalLock_KEY
		port map (
			clk      => clk_clk,                                        --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,   --               reset.reset_n
			address  => key_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => key_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => key_external_export                             -- external_connection.export
		);

	sw : component DigitalLock_SW
		port map (
			clk      => clk_clk,                                       --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,  --               reset.reset_n
			address  => sw_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => sw_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => sw_external_export                             -- external_connection.export
		);

	timer : component DigitalLock_TIMER
		port map (
			clk        => clk_clk,                                                 --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,            -- reset.reset_n
			address    => timer_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                                 --   irq.irq
		);

	sysid : component DigitalLock_sysid
		port map (
			clock    => clk_clk,                                                       --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,                  --         reset.reset_n
			readdata => sysid_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => sysid_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	cpu_instruction_master_translator : component digitallock_cpu_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 15,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 15,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                                   --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                            --                     reset.reset
			uav_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => cpu_instruction_master_read,                                               --                          .read
			av_readdata              => cpu_instruction_master_readdata,                                           --                          .readdata
			av_burstcount            => "1",                                                                       --               (terminated)
			av_byteenable            => "1111",                                                                    --               (terminated)
			av_beginbursttransfer    => '0',                                                                       --               (terminated)
			av_begintransfer         => '0',                                                                       --               (terminated)
			av_chipselect            => '0',                                                                       --               (terminated)
			av_readdatavalid         => open,                                                                      --               (terminated)
			av_write                 => '0',                                                                       --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                        --               (terminated)
			av_lock                  => '0',                                                                       --               (terminated)
			av_debugaccess           => '0',                                                                       --               (terminated)
			uav_clken                => open,                                                                      --               (terminated)
			av_clken                 => '1',                                                                       --               (terminated)
			uav_response             => "00",                                                                      --               (terminated)
			av_response              => open,                                                                      --               (terminated)
			uav_writeresponserequest => open,                                                                      --               (terminated)
			uav_writeresponsevalid   => '0',                                                                       --               (terminated)
			av_writeresponserequest  => '0',                                                                       --               (terminated)
			av_writeresponsevalid    => open                                                                       --               (terminated)
		);

	cpu_data_master_translator : component digitallock_cpu_data_master_translator
		generic map (
			AV_ADDRESS_W                => 15,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 15,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 1
		)
		port map (
			clk                      => clk_clk,                                                            --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                     --                     reset.reset
			uav_address              => cpu_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => cpu_data_master_byteenable,                                         --                          .byteenable
			av_read                  => cpu_data_master_read,                                               --                          .read
			av_readdata              => cpu_data_master_readdata,                                           --                          .readdata
			av_write                 => cpu_data_master_write,                                              --                          .write
			av_writedata             => cpu_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => cpu_data_master_debugaccess,                                        --                          .debugaccess
			av_burstcount            => "1",                                                                --               (terminated)
			av_beginbursttransfer    => '0',                                                                --               (terminated)
			av_begintransfer         => '0',                                                                --               (terminated)
			av_chipselect            => '0',                                                                --               (terminated)
			av_readdatavalid         => open,                                                               --               (terminated)
			av_lock                  => '0',                                                                --               (terminated)
			uav_clken                => open,                                                               --               (terminated)
			av_clken                 => '1',                                                                --               (terminated)
			uav_response             => "00",                                                               --               (terminated)
			av_response              => open,                                                               --               (terminated)
			uav_writeresponserequest => open,                                                               --               (terminated)
			uav_writeresponsevalid   => '0',                                                                --               (terminated)
			av_writeresponserequest  => '0',                                                                --               (terminated)
			av_writeresponsevalid    => open                                                                --               (terminated)
		);

	cpu_jtag_debug_module_translator : component digitallock_cpu_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 15,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                   --                    reset.reset
			uav_address              => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                             --              (terminated)
			av_burstcount            => open,                                                                             --              (terminated)
			av_readdatavalid         => '0',                                                                              --              (terminated)
			av_writebyteenable       => open,                                                                             --              (terminated)
			av_lock                  => open,                                                                             --              (terminated)
			av_chipselect            => open,                                                                             --              (terminated)
			av_clken                 => open,                                                                             --              (terminated)
			uav_clken                => '0',                                                                              --              (terminated)
			av_outputenable          => open,                                                                             --              (terminated)
			uav_response             => open,                                                                             --              (terminated)
			av_response              => "00",                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                               --              (terminated)
		);

	in_ram_s1_translator : component digitallock_in_ram_s1_translator
		generic map (
			AV_ADDRESS_W                   => 11,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 15,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                              --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                   --                    reset.reset
			uav_address              => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => in_ram_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => in_ram_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => in_ram_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => in_ram_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => in_ram_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => in_ram_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_clken                 => in_ram_s1_translator_avalon_anti_slave_0_clken,                       --                         .clken
			av_read                  => open,                                                                 --              (terminated)
			av_begintransfer         => open,                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                 --              (terminated)
			av_burstcount            => open,                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                 --              (terminated)
			av_lock                  => open,                                                                 --              (terminated)
			uav_clken                => '0',                                                                  --              (terminated)
			av_debugaccess           => open,                                                                 --              (terminated)
			av_outputenable          => open,                                                                 --              (terminated)
			uav_response             => open,                                                                 --              (terminated)
			av_response              => "00",                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                   --              (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator : component digitallock_jtag_uart_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 15,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                     --                    reset.reset
			uav_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                   --              (terminated)
			av_burstcount            => open,                                                                                   --              (terminated)
			av_byteenable            => open,                                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                   --              (terminated)
			av_lock                  => open,                                                                                   --              (terminated)
			av_clken                 => open,                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                    --              (terminated)
			av_debugaccess           => open,                                                                                   --              (terminated)
			av_outputenable          => open,                                                                                   --              (terminated)
			uav_response             => open,                                                                                   --              (terminated)
			av_response              => "00",                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                     --              (terminated)
		);

	hex_s1_translator : component digitallock_hex_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 15,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                           --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                --                    reset.reset
			uav_address              => hex_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => hex_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => hex_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => hex_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => hex_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => hex_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => hex_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => hex_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => hex_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => hex_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => hex_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => hex_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => hex_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => hex_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => hex_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => hex_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                              --              (terminated)
			av_begintransfer         => open,                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                              --              (terminated)
			av_burstcount            => open,                                                              --              (terminated)
			av_byteenable            => open,                                                              --              (terminated)
			av_readdatavalid         => '0',                                                               --              (terminated)
			av_waitrequest           => '0',                                                               --              (terminated)
			av_writebyteenable       => open,                                                              --              (terminated)
			av_lock                  => open,                                                              --              (terminated)
			av_clken                 => open,                                                              --              (terminated)
			uav_clken                => '0',                                                               --              (terminated)
			av_debugaccess           => open,                                                              --              (terminated)
			av_outputenable          => open,                                                              --              (terminated)
			uav_response             => open,                                                              --              (terminated)
			av_response              => "00",                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                              --              (terminated)
			av_writeresponserequest  => open,                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                --              (terminated)
		);

	ledg_s1_translator : component digitallock_hex_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 15,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                            --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                 --                    reset.reset
			uav_address              => ledg_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => ledg_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => ledg_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => ledg_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => ledg_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => ledg_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => ledg_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => ledg_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                               --              (terminated)
			av_begintransfer         => open,                                                               --              (terminated)
			av_beginbursttransfer    => open,                                                               --              (terminated)
			av_burstcount            => open,                                                               --              (terminated)
			av_byteenable            => open,                                                               --              (terminated)
			av_readdatavalid         => '0',                                                                --              (terminated)
			av_waitrequest           => '0',                                                                --              (terminated)
			av_writebyteenable       => open,                                                               --              (terminated)
			av_lock                  => open,                                                               --              (terminated)
			av_clken                 => open,                                                               --              (terminated)
			uav_clken                => '0',                                                                --              (terminated)
			av_debugaccess           => open,                                                               --              (terminated)
			av_outputenable          => open,                                                               --              (terminated)
			uav_response             => open,                                                               --              (terminated)
			av_response              => "00",                                                               --              (terminated)
			uav_writeresponserequest => '0',                                                                --              (terminated)
			uav_writeresponsevalid   => open,                                                               --              (terminated)
			av_writeresponserequest  => open,                                                               --              (terminated)
			av_writeresponsevalid    => '0'                                                                 --              (terminated)
		);

	ledr_s1_translator : component digitallock_hex_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 15,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                            --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                 --                    reset.reset
			uav_address              => ledr_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => ledr_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => ledr_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => ledr_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => ledr_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => ledr_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => ledr_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => ledr_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                               --              (terminated)
			av_begintransfer         => open,                                                               --              (terminated)
			av_beginbursttransfer    => open,                                                               --              (terminated)
			av_burstcount            => open,                                                               --              (terminated)
			av_byteenable            => open,                                                               --              (terminated)
			av_readdatavalid         => '0',                                                                --              (terminated)
			av_waitrequest           => '0',                                                                --              (terminated)
			av_writebyteenable       => open,                                                               --              (terminated)
			av_lock                  => open,                                                               --              (terminated)
			av_clken                 => open,                                                               --              (terminated)
			uav_clken                => '0',                                                                --              (terminated)
			av_debugaccess           => open,                                                               --              (terminated)
			av_outputenable          => open,                                                               --              (terminated)
			uav_response             => open,                                                               --              (terminated)
			av_response              => "00",                                                               --              (terminated)
			uav_writeresponserequest => '0',                                                                --              (terminated)
			uav_writeresponsevalid   => open,                                                               --              (terminated)
			av_writeresponserequest  => open,                                                               --              (terminated)
			av_writeresponsevalid    => '0'                                                                 --              (terminated)
		);

	key_s1_translator : component digitallock_key_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 15,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                           --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                --                    reset.reset
			uav_address              => key_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => key_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => key_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => key_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => key_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => key_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => key_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => key_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                              --              (terminated)
			av_read                  => open,                                                              --              (terminated)
			av_writedata             => open,                                                              --              (terminated)
			av_begintransfer         => open,                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                              --              (terminated)
			av_burstcount            => open,                                                              --              (terminated)
			av_byteenable            => open,                                                              --              (terminated)
			av_readdatavalid         => '0',                                                               --              (terminated)
			av_waitrequest           => '0',                                                               --              (terminated)
			av_writebyteenable       => open,                                                              --              (terminated)
			av_lock                  => open,                                                              --              (terminated)
			av_chipselect            => open,                                                              --              (terminated)
			av_clken                 => open,                                                              --              (terminated)
			uav_clken                => '0',                                                               --              (terminated)
			av_debugaccess           => open,                                                              --              (terminated)
			av_outputenable          => open,                                                              --              (terminated)
			uav_response             => open,                                                              --              (terminated)
			av_response              => "00",                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                              --              (terminated)
			av_writeresponserequest  => open,                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                --              (terminated)
		);

	sw_s1_translator : component digitallock_key_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 15,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                          --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                               --                    reset.reset
			uav_address              => sw_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sw_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sw_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sw_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sw_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => sw_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                             --              (terminated)
			av_read                  => open,                                                             --              (terminated)
			av_writedata             => open,                                                             --              (terminated)
			av_begintransfer         => open,                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                             --              (terminated)
			av_burstcount            => open,                                                             --              (terminated)
			av_byteenable            => open,                                                             --              (terminated)
			av_readdatavalid         => '0',                                                              --              (terminated)
			av_waitrequest           => '0',                                                              --              (terminated)
			av_writebyteenable       => open,                                                             --              (terminated)
			av_lock                  => open,                                                             --              (terminated)
			av_chipselect            => open,                                                             --              (terminated)
			av_clken                 => open,                                                             --              (terminated)
			uav_clken                => '0',                                                              --              (terminated)
			av_debugaccess           => open,                                                             --              (terminated)
			av_outputenable          => open,                                                             --              (terminated)
			uav_response             => open,                                                             --              (terminated)
			av_response              => "00",                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                             --              (terminated)
			av_writeresponserequest  => open,                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                               --              (terminated)
		);

	timer_s1_translator : component digitallock_timer_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 15,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                             --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                  --                    reset.reset
			uav_address              => timer_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => timer_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => timer_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => timer_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => timer_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => timer_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => timer_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => timer_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => timer_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                --              (terminated)
			av_begintransfer         => open,                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                --              (terminated)
			av_burstcount            => open,                                                                --              (terminated)
			av_byteenable            => open,                                                                --              (terminated)
			av_readdatavalid         => '0',                                                                 --              (terminated)
			av_waitrequest           => '0',                                                                 --              (terminated)
			av_writebyteenable       => open,                                                                --              (terminated)
			av_lock                  => open,                                                                --              (terminated)
			av_clken                 => open,                                                                --              (terminated)
			uav_clken                => '0',                                                                 --              (terminated)
			av_debugaccess           => open,                                                                --              (terminated)
			av_outputenable          => open,                                                                --              (terminated)
			uav_response             => open,                                                                --              (terminated)
			av_response              => "00",                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                  --              (terminated)
		);

	sysid_control_slave_translator : component digitallock_sysid_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 15,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                        --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                             --                    reset.reset
			uav_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sysid_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => sysid_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                           --              (terminated)
			av_read                  => open,                                                                           --              (terminated)
			av_writedata             => open,                                                                           --              (terminated)
			av_begintransfer         => open,                                                                           --              (terminated)
			av_beginbursttransfer    => open,                                                                           --              (terminated)
			av_burstcount            => open,                                                                           --              (terminated)
			av_byteenable            => open,                                                                           --              (terminated)
			av_readdatavalid         => '0',                                                                            --              (terminated)
			av_waitrequest           => '0',                                                                            --              (terminated)
			av_writebyteenable       => open,                                                                           --              (terminated)
			av_lock                  => open,                                                                           --              (terminated)
			av_chipselect            => open,                                                                           --              (terminated)
			av_clken                 => open,                                                                           --              (terminated)
			uav_clken                => '0',                                                                            --              (terminated)
			av_debugaccess           => open,                                                                           --              (terminated)
			av_outputenable          => open,                                                                           --              (terminated)
			uav_response             => open,                                                                           --              (terminated)
			av_response              => "00",                                                                           --              (terminated)
			uav_writeresponserequest => '0',                                                                            --              (terminated)
			uav_writeresponsevalid   => open,                                                                           --              (terminated)
			av_writeresponserequest  => open,                                                                           --              (terminated)
			av_writeresponsevalid    => '0'                                                                             --              (terminated)
		);

	cpu_instruction_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 83,
			PKT_PROTECTION_L          => 81,
			PKT_BEGIN_BURST           => 70,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			PKT_BURST_TYPE_H          => 67,
			PKT_BURST_TYPE_L          => 66,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 57,
			PKT_ADDR_H                => 50,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 51,
			PKT_TRANS_POSTED          => 52,
			PKT_TRANS_WRITE           => 53,
			PKT_TRANS_READ            => 54,
			PKT_TRANS_LOCK            => 55,
			PKT_TRANS_EXCLUSIVE       => 56,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 79,
			PKT_DEST_ID_L             => 76,
			PKT_THREAD_ID_H           => 80,
			PKT_THREAD_ID_L           => 80,
			PKT_CACHE_H               => 87,
			PKT_CACHE_L               => 84,
			PKT_DATA_SIDEBAND_H       => 69,
			PKT_DATA_SIDEBAND_L       => 69,
			PKT_QOS_H                 => 71,
			PKT_QOS_L                 => 71,
			PKT_ADDR_SIDEBAND_H       => 68,
			PKT_ADDR_SIDEBAND_L       => 68,
			PKT_RESPONSE_STATUS_H     => 89,
			PKT_RESPONSE_STATUS_L     => 88,
			ST_DATA_W                 => 90,
			ST_CHANNEL_W              => 10,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                            --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			av_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_src_valid,                                                             --        rp.valid
			rp_data                 => rsp_xbar_mux_src_data,                                                              --          .data
			rp_channel              => rsp_xbar_mux_src_channel,                                                           --          .channel
			rp_startofpacket        => rsp_xbar_mux_src_startofpacket,                                                     --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_src_endofpacket,                                                       --          .endofpacket
			rp_ready                => rsp_xbar_mux_src_ready,                                                             --          .ready
			av_response             => open,                                                                               -- (terminated)
			av_writeresponserequest => '0',                                                                                -- (terminated)
			av_writeresponsevalid   => open                                                                                -- (terminated)
		);

	cpu_data_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 83,
			PKT_PROTECTION_L          => 81,
			PKT_BEGIN_BURST           => 70,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			PKT_BURST_TYPE_H          => 67,
			PKT_BURST_TYPE_L          => 66,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 57,
			PKT_ADDR_H                => 50,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 51,
			PKT_TRANS_POSTED          => 52,
			PKT_TRANS_WRITE           => 53,
			PKT_TRANS_READ            => 54,
			PKT_TRANS_LOCK            => 55,
			PKT_TRANS_EXCLUSIVE       => 56,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 79,
			PKT_DEST_ID_L             => 76,
			PKT_THREAD_ID_H           => 80,
			PKT_THREAD_ID_L           => 80,
			PKT_CACHE_H               => 87,
			PKT_CACHE_L               => 84,
			PKT_DATA_SIDEBAND_H       => 69,
			PKT_DATA_SIDEBAND_L       => 69,
			PKT_QOS_H                 => 71,
			PKT_QOS_L                 => 71,
			PKT_ADDR_SIDEBAND_H       => 68,
			PKT_ADDR_SIDEBAND_L       => 68,
			PKT_RESPONSE_STATUS_H     => 89,
			PKT_RESPONSE_STATUS_L     => 88,
			ST_DATA_W                 => 90,
			ST_CHANNEL_W              => 10,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                     --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			av_address              => cpu_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_001_src_valid,                                                  --        rp.valid
			rp_data                 => rsp_xbar_mux_001_src_data,                                                   --          .data
			rp_channel              => rsp_xbar_mux_001_src_channel,                                                --          .channel
			rp_startofpacket        => rsp_xbar_mux_001_src_startofpacket,                                          --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_001_src_endofpacket,                                            --          .endofpacket
			rp_ready                => rsp_xbar_mux_001_src_ready,                                                  --          .ready
			av_response             => open,                                                                        -- (terminated)
			av_writeresponserequest => '0',                                                                         -- (terminated)
			av_writeresponsevalid   => open                                                                         -- (terminated)
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 50,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 51,
			PKT_TRANS_POSTED          => 52,
			PKT_TRANS_WRITE           => 53,
			PKT_TRANS_READ            => 54,
			PKT_TRANS_LOCK            => 55,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 79,
			PKT_DEST_ID_L             => 76,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 57,
			PKT_PROTECTION_H          => 83,
			PKT_PROTECTION_L          => 81,
			PKT_RESPONSE_STATUS_H     => 89,
			PKT_RESPONSE_STATUS_L     => 88,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 90,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                             --       clk_reset.reset
			m0_address              => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                     --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                     --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                      --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                               --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                   --                .channel
			rf_sink_ready           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                         --     (terminated)
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 91,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                             -- clk_reset.reset
			in_data           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                       -- (terminated)
			csr_read          => '0',                                                                                        -- (terminated)
			csr_write         => '0',                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                         -- (terminated)
			almost_full_data  => open,                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                       -- (terminated)
			in_empty          => '0',                                                                                        -- (terminated)
			out_empty         => open,                                                                                       -- (terminated)
			in_error          => '0',                                                                                        -- (terminated)
			out_error         => open,                                                                                       -- (terminated)
			in_channel        => '0',                                                                                        -- (terminated)
			out_channel       => open                                                                                        -- (terminated)
		);

	in_ram_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 50,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 51,
			PKT_TRANS_POSTED          => 52,
			PKT_TRANS_WRITE           => 53,
			PKT_TRANS_READ            => 54,
			PKT_TRANS_LOCK            => 55,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 79,
			PKT_DEST_ID_L             => 76,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 57,
			PKT_PROTECTION_H          => 83,
			PKT_PROTECTION_L          => 81,
			PKT_RESPONSE_STATUS_H     => 89,
			PKT_RESPONSE_STATUS_L     => 88,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 90,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                        --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                             --       clk_reset.reset
			m0_address              => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => in_ram_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => in_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => in_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => in_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => in_ram_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => in_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_001_src_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_mux_001_src_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_mux_001_src_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_mux_001_src_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_001_src_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_mux_001_src_channel,                                                   --                .channel
			rf_sink_ready           => in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => in_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => in_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => in_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => in_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => in_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => in_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                             --     (terminated)
		);

	in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 91,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                        --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			in_data           => in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => in_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => in_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 50,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 51,
			PKT_TRANS_POSTED          => 52,
			PKT_TRANS_WRITE           => 53,
			PKT_TRANS_READ            => 54,
			PKT_TRANS_LOCK            => 55,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 79,
			PKT_DEST_ID_L             => 76,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 57,
			PKT_PROTECTION_H          => 83,
			PKT_PROTECTION_L          => 81,
			PKT_RESPONSE_STATUS_H     => 89,
			PKT_RESPONSE_STATUS_L     => 88,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 90,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                          --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                               --       clk_reset.reset
			m0_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src2_ready,                                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src2_valid,                                                                    --                .valid
			cp_data                 => cmd_xbar_demux_001_src2_data,                                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src2_startofpacket,                                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src2_endofpacket,                                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src2_channel,                                                                  --                .channel
			rf_sink_ready           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                               --     (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 91,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                          --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                               -- clk_reset.reset
			in_data           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                             -- (terminated)
			csr_read          => '0',                                                                                              -- (terminated)
			csr_write         => '0',                                                                                              -- (terminated)
			csr_readdata      => open,                                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                               -- (terminated)
			almost_full_data  => open,                                                                                             -- (terminated)
			almost_empty_data => open,                                                                                             -- (terminated)
			in_empty          => '0',                                                                                              -- (terminated)
			out_empty         => open,                                                                                             -- (terminated)
			in_error          => '0',                                                                                              -- (terminated)
			out_error         => open,                                                                                             -- (terminated)
			in_channel        => '0',                                                                                              -- (terminated)
			out_channel       => open                                                                                              -- (terminated)
		);

	hex_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 50,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 51,
			PKT_TRANS_POSTED          => 52,
			PKT_TRANS_WRITE           => 53,
			PKT_TRANS_READ            => 54,
			PKT_TRANS_LOCK            => 55,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 79,
			PKT_DEST_ID_L             => 76,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 57,
			PKT_PROTECTION_H          => 83,
			PKT_PROTECTION_L          => 81,
			PKT_RESPONSE_STATUS_H     => 89,
			PKT_RESPONSE_STATUS_L     => 88,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 90,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                     --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                          --       clk_reset.reset
			m0_address              => hex_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => hex_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => hex_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => hex_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => hex_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => hex_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => hex_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => hex_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => hex_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => hex_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => hex_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => hex_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => hex_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => hex_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => hex_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => hex_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src3_ready,                                               --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src3_valid,                                               --                .valid
			cp_data                 => cmd_xbar_demux_001_src3_data,                                                --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src3_startofpacket,                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src3_endofpacket,                                         --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src3_channel,                                             --                .channel
			rf_sink_ready           => hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => hex_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => hex_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => hex_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => hex_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => hex_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => hex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => hex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => hex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => hex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => hex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => hex_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                          --     (terminated)
		);

	hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 91,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                          -- clk_reset.reset
			in_data           => hex_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => hex_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => hex_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => hex_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => hex_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => hex_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                        -- (terminated)
			csr_read          => '0',                                                                         -- (terminated)
			csr_write         => '0',                                                                         -- (terminated)
			csr_readdata      => open,                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                          -- (terminated)
			almost_full_data  => open,                                                                        -- (terminated)
			almost_empty_data => open,                                                                        -- (terminated)
			in_empty          => '0',                                                                         -- (terminated)
			out_empty         => open,                                                                        -- (terminated)
			in_error          => '0',                                                                         -- (terminated)
			out_error         => open,                                                                        -- (terminated)
			in_channel        => '0',                                                                         -- (terminated)
			out_channel       => open                                                                         -- (terminated)
		);

	ledg_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 50,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 51,
			PKT_TRANS_POSTED          => 52,
			PKT_TRANS_WRITE           => 53,
			PKT_TRANS_READ            => 54,
			PKT_TRANS_LOCK            => 55,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 79,
			PKT_DEST_ID_L             => 76,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 57,
			PKT_PROTECTION_H          => 83,
			PKT_PROTECTION_L          => 81,
			PKT_RESPONSE_STATUS_H     => 89,
			PKT_RESPONSE_STATUS_L     => 88,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 90,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                      --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                           --       clk_reset.reset
			m0_address              => ledg_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => ledg_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => ledg_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => ledg_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src4_ready,                                                --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src4_valid,                                                --                .valid
			cp_data                 => cmd_xbar_demux_001_src4_data,                                                 --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src4_startofpacket,                                        --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src4_endofpacket,                                          --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src4_channel,                                              --                .channel
			rf_sink_ready           => ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                         --     (terminated)
			m0_writeresponserequest => open,                                                                         --     (terminated)
			m0_writeresponsevalid   => '0'                                                                           --     (terminated)
		);

	ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 91,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                      --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                           -- clk_reset.reset
			in_data           => ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                         -- (terminated)
			csr_read          => '0',                                                                          -- (terminated)
			csr_write         => '0',                                                                          -- (terminated)
			csr_readdata      => open,                                                                         -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                           -- (terminated)
			almost_full_data  => open,                                                                         -- (terminated)
			almost_empty_data => open,                                                                         -- (terminated)
			in_empty          => '0',                                                                          -- (terminated)
			out_empty         => open,                                                                         -- (terminated)
			in_error          => '0',                                                                          -- (terminated)
			out_error         => open,                                                                         -- (terminated)
			in_channel        => '0',                                                                          -- (terminated)
			out_channel       => open                                                                          -- (terminated)
		);

	ledr_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 50,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 51,
			PKT_TRANS_POSTED          => 52,
			PKT_TRANS_WRITE           => 53,
			PKT_TRANS_READ            => 54,
			PKT_TRANS_LOCK            => 55,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 79,
			PKT_DEST_ID_L             => 76,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 57,
			PKT_PROTECTION_H          => 83,
			PKT_PROTECTION_L          => 81,
			PKT_RESPONSE_STATUS_H     => 89,
			PKT_RESPONSE_STATUS_L     => 88,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 90,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                      --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                           --       clk_reset.reset
			m0_address              => ledr_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => ledr_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => ledr_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => ledr_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src5_ready,                                                --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src5_valid,                                                --                .valid
			cp_data                 => cmd_xbar_demux_001_src5_data,                                                 --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src5_startofpacket,                                        --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src5_endofpacket,                                          --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src5_channel,                                              --                .channel
			rf_sink_ready           => ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                         --     (terminated)
			m0_writeresponserequest => open,                                                                         --     (terminated)
			m0_writeresponsevalid   => '0'                                                                           --     (terminated)
		);

	ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 91,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                      --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                           -- clk_reset.reset
			in_data           => ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                         -- (terminated)
			csr_read          => '0',                                                                          -- (terminated)
			csr_write         => '0',                                                                          -- (terminated)
			csr_readdata      => open,                                                                         -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                           -- (terminated)
			almost_full_data  => open,                                                                         -- (terminated)
			almost_empty_data => open,                                                                         -- (terminated)
			in_empty          => '0',                                                                          -- (terminated)
			out_empty         => open,                                                                         -- (terminated)
			in_error          => '0',                                                                          -- (terminated)
			out_error         => open,                                                                         -- (terminated)
			in_channel        => '0',                                                                          -- (terminated)
			out_channel       => open                                                                          -- (terminated)
		);

	key_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 50,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 51,
			PKT_TRANS_POSTED          => 52,
			PKT_TRANS_WRITE           => 53,
			PKT_TRANS_READ            => 54,
			PKT_TRANS_LOCK            => 55,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 79,
			PKT_DEST_ID_L             => 76,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 57,
			PKT_PROTECTION_H          => 83,
			PKT_PROTECTION_L          => 81,
			PKT_RESPONSE_STATUS_H     => 89,
			PKT_RESPONSE_STATUS_L     => 88,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 90,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                     --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                          --       clk_reset.reset
			m0_address              => key_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => key_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => key_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => key_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => key_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => key_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => key_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => key_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => key_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src6_ready,                                               --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src6_valid,                                               --                .valid
			cp_data                 => cmd_xbar_demux_001_src6_data,                                                --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src6_startofpacket,                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src6_endofpacket,                                         --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src6_channel,                                             --                .channel
			rf_sink_ready           => key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => key_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                          --     (terminated)
		);

	key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 91,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                          -- clk_reset.reset
			in_data           => key_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                        -- (terminated)
			csr_read          => '0',                                                                         -- (terminated)
			csr_write         => '0',                                                                         -- (terminated)
			csr_readdata      => open,                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                          -- (terminated)
			almost_full_data  => open,                                                                        -- (terminated)
			almost_empty_data => open,                                                                        -- (terminated)
			in_empty          => '0',                                                                         -- (terminated)
			out_empty         => open,                                                                        -- (terminated)
			in_error          => '0',                                                                         -- (terminated)
			out_error         => open,                                                                        -- (terminated)
			in_channel        => '0',                                                                         -- (terminated)
			out_channel       => open                                                                         -- (terminated)
		);

	sw_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 50,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 51,
			PKT_TRANS_POSTED          => 52,
			PKT_TRANS_WRITE           => 53,
			PKT_TRANS_READ            => 54,
			PKT_TRANS_LOCK            => 55,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 79,
			PKT_DEST_ID_L             => 76,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 57,
			PKT_PROTECTION_H          => 83,
			PKT_PROTECTION_L          => 81,
			PKT_RESPONSE_STATUS_H     => 89,
			PKT_RESPONSE_STATUS_L     => 88,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 90,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                    --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                         --       clk_reset.reset
			m0_address              => sw_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sw_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sw_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sw_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sw_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sw_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sw_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src7_ready,                                              --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src7_valid,                                              --                .valid
			cp_data                 => cmd_xbar_demux_001_src7_data,                                               --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src7_startofpacket,                                      --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src7_endofpacket,                                        --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src7_channel,                                            --                .channel
			rf_sink_ready           => sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                         --     (terminated)
		);

	sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 91,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                    --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                         -- clk_reset.reset
			in_data           => sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                       -- (terminated)
			csr_read          => '0',                                                                        -- (terminated)
			csr_write         => '0',                                                                        -- (terminated)
			csr_readdata      => open,                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                         -- (terminated)
			almost_full_data  => open,                                                                       -- (terminated)
			almost_empty_data => open,                                                                       -- (terminated)
			in_empty          => '0',                                                                        -- (terminated)
			out_empty         => open,                                                                       -- (terminated)
			in_error          => '0',                                                                        -- (terminated)
			out_error         => open,                                                                       -- (terminated)
			in_channel        => '0',                                                                        -- (terminated)
			out_channel       => open                                                                        -- (terminated)
		);

	timer_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 50,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 51,
			PKT_TRANS_POSTED          => 52,
			PKT_TRANS_WRITE           => 53,
			PKT_TRANS_READ            => 54,
			PKT_TRANS_LOCK            => 55,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 79,
			PKT_DEST_ID_L             => 76,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 57,
			PKT_PROTECTION_H          => 83,
			PKT_PROTECTION_L          => 81,
			PKT_RESPONSE_STATUS_H     => 89,
			PKT_RESPONSE_STATUS_L     => 88,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 90,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                       --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                            --       clk_reset.reset
			m0_address              => timer_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src8_ready,                                                 --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src8_valid,                                                 --                .valid
			cp_data                 => cmd_xbar_demux_001_src8_data,                                                  --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src8_startofpacket,                                         --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src8_endofpacket,                                           --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src8_channel,                                               --                .channel
			rf_sink_ready           => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                            --     (terminated)
		);

	timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 91,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                       --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                            -- clk_reset.reset
			in_data           => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                          -- (terminated)
			csr_read          => '0',                                                                           -- (terminated)
			csr_write         => '0',                                                                           -- (terminated)
			csr_readdata      => open,                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                            -- (terminated)
			almost_full_data  => open,                                                                          -- (terminated)
			almost_empty_data => open,                                                                          -- (terminated)
			in_empty          => '0',                                                                           -- (terminated)
			out_empty         => open,                                                                          -- (terminated)
			in_error          => '0',                                                                           -- (terminated)
			out_error         => open,                                                                          -- (terminated)
			in_channel        => '0',                                                                           -- (terminated)
			out_channel       => open                                                                           -- (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 50,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 51,
			PKT_TRANS_POSTED          => 52,
			PKT_TRANS_WRITE           => 53,
			PKT_TRANS_READ            => 54,
			PKT_TRANS_LOCK            => 55,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 79,
			PKT_DEST_ID_L             => 76,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 57,
			PKT_PROTECTION_H          => 83,
			PKT_PROTECTION_L          => 81,
			PKT_RESPONSE_STATUS_H     => 89,
			PKT_RESPONSE_STATUS_L     => 88,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 90,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                  --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                       --       clk_reset.reset
			m0_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src9_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src9_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_demux_001_src9_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src9_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src9_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src9_channel,                                                          --                .channel
			rf_sink_ready           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                     --     (terminated)
			m0_writeresponserequest => open,                                                                                     --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                       --     (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 91,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                  --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                       -- clk_reset.reset
			in_data           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                     -- (terminated)
			csr_read          => '0',                                                                                      -- (terminated)
			csr_write         => '0',                                                                                      -- (terminated)
			csr_readdata      => open,                                                                                     -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                       -- (terminated)
			almost_full_data  => open,                                                                                     -- (terminated)
			almost_empty_data => open,                                                                                     -- (terminated)
			in_empty          => '0',                                                                                      -- (terminated)
			out_empty         => open,                                                                                     -- (terminated)
			in_error          => '0',                                                                                      -- (terminated)
			out_error         => open,                                                                                     -- (terminated)
			in_channel        => '0',                                                                                      -- (terminated)
			out_channel       => open                                                                                      -- (terminated)
		);

	addr_router : component DigitalLock_addr_router
		port map (
			sink_ready         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                              --       src.ready
			src_valid          => addr_router_src_valid,                                                              --          .valid
			src_data           => addr_router_src_data,                                                               --          .data
			src_channel        => addr_router_src_channel,                                                            --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                         --          .endofpacket
		);

	addr_router_001 : component DigitalLock_addr_router_001
		port map (
			sink_ready         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                   --       src.ready
			src_valid          => addr_router_001_src_valid,                                                   --          .valid
			src_data           => addr_router_001_src_data,                                                    --          .data
			src_channel        => addr_router_001_src_channel,                                                 --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                           --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                              --          .endofpacket
		);

	id_router : component DigitalLock_id_router
		port map (
			sink_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                              --       src.ready
			src_valid          => id_router_src_valid,                                                              --          .valid
			src_data           => id_router_src_data,                                                               --          .data
			src_channel        => id_router_src_channel,                                                            --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                         --          .endofpacket
		);

	id_router_001 : component DigitalLock_id_router
		port map (
			sink_ready         => in_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => in_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => in_ram_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => in_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => in_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                              --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                   -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                              --       src.ready
			src_valid          => id_router_001_src_valid,                                              --          .valid
			src_data           => id_router_001_src_data,                                               --          .data
			src_channel        => id_router_001_src_channel,                                            --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                         --          .endofpacket
		);

	id_router_002 : component DigitalLock_id_router_002
		port map (
			sink_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                                --       src.ready
			src_valid          => id_router_002_src_valid,                                                                --          .valid
			src_data           => id_router_002_src_data,                                                                 --          .data
			src_channel        => id_router_002_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                           --          .endofpacket
		);

	id_router_003 : component DigitalLock_id_router_002
		port map (
			sink_ready         => hex_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => hex_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => hex_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => hex_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => hex_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                           --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                           --       src.ready
			src_valid          => id_router_003_src_valid,                                           --          .valid
			src_data           => id_router_003_src_data,                                            --          .data
			src_channel        => id_router_003_src_channel,                                         --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                   --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                      --          .endofpacket
		);

	id_router_004 : component DigitalLock_id_router_002
		port map (
			sink_ready         => ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => ledg_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                            --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                 -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                            --       src.ready
			src_valid          => id_router_004_src_valid,                                            --          .valid
			src_data           => id_router_004_src_data,                                             --          .data
			src_channel        => id_router_004_src_channel,                                          --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                    --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                       --          .endofpacket
		);

	id_router_005 : component DigitalLock_id_router_002
		port map (
			sink_ready         => ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => ledr_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                            --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                 -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                            --       src.ready
			src_valid          => id_router_005_src_valid,                                            --          .valid
			src_data           => id_router_005_src_data,                                             --          .data
			src_channel        => id_router_005_src_channel,                                          --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                    --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                       --          .endofpacket
		);

	id_router_006 : component DigitalLock_id_router_002
		port map (
			sink_ready         => key_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => key_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => key_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                           --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                           --       src.ready
			src_valid          => id_router_006_src_valid,                                           --          .valid
			src_data           => id_router_006_src_data,                                            --          .data
			src_channel        => id_router_006_src_channel,                                         --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                   --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                      --          .endofpacket
		);

	id_router_007 : component DigitalLock_id_router_002
		port map (
			sink_ready         => sw_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sw_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sw_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                          --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                               -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                          --       src.ready
			src_valid          => id_router_007_src_valid,                                          --          .valid
			src_data           => id_router_007_src_data,                                           --          .data
			src_channel        => id_router_007_src_channel,                                        --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                  --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                     --          .endofpacket
		);

	id_router_008 : component DigitalLock_id_router_002
		port map (
			sink_ready         => timer_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                             --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                  -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                             --       src.ready
			src_valid          => id_router_008_src_valid,                                             --          .valid
			src_data           => id_router_008_src_data,                                              --          .data
			src_channel        => id_router_008_src_channel,                                           --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                     --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                        --          .endofpacket
		);

	id_router_009 : component DigitalLock_id_router_002
		port map (
			sink_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                        --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                                        --       src.ready
			src_valid          => id_router_009_src_valid,                                                        --          .valid
			src_data           => id_router_009_src_data,                                                         --          .data
			src_channel        => id_router_009_src_channel,                                                      --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                                --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                                   --          .endofpacket
		);

	rst_controller : component digitallock_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 2,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => cpu_jtag_debug_module_reset_reset, -- reset_in0.reset
			reset_in1  => cpu_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk        => clk_clk,                           --       clk.clk
			reset_out  => rst_controller_reset_out_reset,    -- reset_out.reset
			reset_req  => open,                              -- (terminated)
			reset_in2  => '0',                               -- (terminated)
			reset_in3  => '0',                               -- (terminated)
			reset_in4  => '0',                               -- (terminated)
			reset_in5  => '0',                               -- (terminated)
			reset_in6  => '0',                               -- (terminated)
			reset_in7  => '0',                               -- (terminated)
			reset_in8  => '0',                               -- (terminated)
			reset_in9  => '0',                               -- (terminated)
			reset_in10 => '0',                               -- (terminated)
			reset_in11 => '0',                               -- (terminated)
			reset_in12 => '0',                               -- (terminated)
			reset_in13 => '0',                               -- (terminated)
			reset_in14 => '0',                               -- (terminated)
			reset_in15 => '0'                                -- (terminated)
		);

	rst_controller_001 : component digitallock_rst_controller_001
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 1
		)
		port map (
			reset_in0  => cpu_jtag_debug_module_reset_reset,      -- reset_in0.reset
			clk        => clk_clk,                                --       clk.clk
			reset_out  => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req  => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_in1  => '0',                                    -- (terminated)
			reset_in2  => '0',                                    -- (terminated)
			reset_in3  => '0',                                    -- (terminated)
			reset_in4  => '0',                                    -- (terminated)
			reset_in5  => '0',                                    -- (terminated)
			reset_in6  => '0',                                    -- (terminated)
			reset_in7  => '0',                                    -- (terminated)
			reset_in8  => '0',                                    -- (terminated)
			reset_in9  => '0',                                    -- (terminated)
			reset_in10 => '0',                                    -- (terminated)
			reset_in11 => '0',                                    -- (terminated)
			reset_in12 => '0',                                    -- (terminated)
			reset_in13 => '0',                                    -- (terminated)
			reset_in14 => '0',                                    -- (terminated)
			reset_in15 => '0'                                     -- (terminated)
		);

	cmd_xbar_demux : component DigitalLock_cmd_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_src_ready,             --      sink.ready
			sink_channel       => addr_router_src_channel,           --          .channel
			sink_data          => addr_router_src_data,              --          .data
			sink_startofpacket => addr_router_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_001 : component DigitalLock_cmd_xbar_demux_001
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_001_src_ready,             --      sink.ready
			sink_channel       => addr_router_001_src_channel,           --          .channel
			sink_data          => addr_router_001_src_data,              --          .data
			sink_startofpacket => addr_router_001_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_001_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_001_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_001_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			src2_ready         => cmd_xbar_demux_001_src2_ready,         --      src2.ready
			src2_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			src2_data          => cmd_xbar_demux_001_src2_data,          --          .data
			src2_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			src2_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => cmd_xbar_demux_001_src2_endofpacket,   --          .endofpacket
			src3_ready         => cmd_xbar_demux_001_src3_ready,         --      src3.ready
			src3_valid         => cmd_xbar_demux_001_src3_valid,         --          .valid
			src3_data          => cmd_xbar_demux_001_src3_data,          --          .data
			src3_channel       => cmd_xbar_demux_001_src3_channel,       --          .channel
			src3_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --          .startofpacket
			src3_endofpacket   => cmd_xbar_demux_001_src3_endofpacket,   --          .endofpacket
			src4_ready         => cmd_xbar_demux_001_src4_ready,         --      src4.ready
			src4_valid         => cmd_xbar_demux_001_src4_valid,         --          .valid
			src4_data          => cmd_xbar_demux_001_src4_data,          --          .data
			src4_channel       => cmd_xbar_demux_001_src4_channel,       --          .channel
			src4_startofpacket => cmd_xbar_demux_001_src4_startofpacket, --          .startofpacket
			src4_endofpacket   => cmd_xbar_demux_001_src4_endofpacket,   --          .endofpacket
			src5_ready         => cmd_xbar_demux_001_src5_ready,         --      src5.ready
			src5_valid         => cmd_xbar_demux_001_src5_valid,         --          .valid
			src5_data          => cmd_xbar_demux_001_src5_data,          --          .data
			src5_channel       => cmd_xbar_demux_001_src5_channel,       --          .channel
			src5_startofpacket => cmd_xbar_demux_001_src5_startofpacket, --          .startofpacket
			src5_endofpacket   => cmd_xbar_demux_001_src5_endofpacket,   --          .endofpacket
			src6_ready         => cmd_xbar_demux_001_src6_ready,         --      src6.ready
			src6_valid         => cmd_xbar_demux_001_src6_valid,         --          .valid
			src6_data          => cmd_xbar_demux_001_src6_data,          --          .data
			src6_channel       => cmd_xbar_demux_001_src6_channel,       --          .channel
			src6_startofpacket => cmd_xbar_demux_001_src6_startofpacket, --          .startofpacket
			src6_endofpacket   => cmd_xbar_demux_001_src6_endofpacket,   --          .endofpacket
			src7_ready         => cmd_xbar_demux_001_src7_ready,         --      src7.ready
			src7_valid         => cmd_xbar_demux_001_src7_valid,         --          .valid
			src7_data          => cmd_xbar_demux_001_src7_data,          --          .data
			src7_channel       => cmd_xbar_demux_001_src7_channel,       --          .channel
			src7_startofpacket => cmd_xbar_demux_001_src7_startofpacket, --          .startofpacket
			src7_endofpacket   => cmd_xbar_demux_001_src7_endofpacket,   --          .endofpacket
			src8_ready         => cmd_xbar_demux_001_src8_ready,         --      src8.ready
			src8_valid         => cmd_xbar_demux_001_src8_valid,         --          .valid
			src8_data          => cmd_xbar_demux_001_src8_data,          --          .data
			src8_channel       => cmd_xbar_demux_001_src8_channel,       --          .channel
			src8_startofpacket => cmd_xbar_demux_001_src8_startofpacket, --          .startofpacket
			src8_endofpacket   => cmd_xbar_demux_001_src8_endofpacket,   --          .endofpacket
			src9_ready         => cmd_xbar_demux_001_src9_ready,         --      src9.ready
			src9_valid         => cmd_xbar_demux_001_src9_valid,         --          .valid
			src9_data          => cmd_xbar_demux_001_src9_data,          --          .data
			src9_channel       => cmd_xbar_demux_001_src9_channel,       --          .channel
			src9_startofpacket => cmd_xbar_demux_001_src9_startofpacket, --          .startofpacket
			src9_endofpacket   => cmd_xbar_demux_001_src9_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component DigitalLock_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component DigitalLock_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component DigitalLock_cmd_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component DigitalLock_cmd_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component DigitalLock_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component DigitalLock_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component DigitalLock_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component DigitalLock_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component DigitalLock_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component DigitalLock_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component DigitalLock_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component DigitalLock_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component DigitalLock_rsp_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component DigitalLock_rsp_xbar_mux_001
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data            => rsp_xbar_mux_001_src_data,             --          .data
			src_channel         => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready         => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink4_ready         => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data          => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink5_ready         => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data          => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket   => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready         => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data          => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket   => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink7_ready         => rsp_xbar_demux_007_src0_ready,         --     sink7.ready
			sink7_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink7_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink7_data          => rsp_xbar_demux_007_src0_data,          --          .data
			sink7_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink7_endofpacket   => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			sink8_ready         => rsp_xbar_demux_008_src0_ready,         --     sink8.ready
			sink8_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			sink8_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			sink8_data          => rsp_xbar_demux_008_src0_data,          --          .data
			sink8_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			sink8_endofpacket   => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			sink9_ready         => rsp_xbar_demux_009_src0_ready,         --     sink9.ready
			sink9_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink9_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink9_data          => rsp_xbar_demux_009_src0_data,          --          .data
			sink9_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink9_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	irq_mapper : component DigitalLock_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_d_irq_irq                   --    sender.irq
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	hex_s1_translator_avalon_anti_slave_0_write_ports_inv <= not hex_s1_translator_avalon_anti_slave_0_write;

	ledg_s1_translator_avalon_anti_slave_0_write_ports_inv <= not ledg_s1_translator_avalon_anti_slave_0_write;

	ledr_s1_translator_avalon_anti_slave_0_write_ports_inv <= not ledr_s1_translator_avalon_anti_slave_0_write;

	timer_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_s1_translator_avalon_anti_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of DigitalLock
